module adapter256c8 (
	input clk,
	input reset,
	input in_vld,
	input [255:0] in_data,
	output rdy_in,
	output vld_out,
	output [7:0] data_out,
	input out_rdy
);
	reg [255:0] temp;
	
endmodule

module adapter8c256 (

);

endmodule
